module hello;
    initial begin
        $display("Hello world\n");
    end
endmodule